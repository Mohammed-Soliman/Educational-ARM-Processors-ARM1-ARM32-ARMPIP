// flip-flop with enable and async reset
module flopenr #(parameter WIDTH = 8) (
input logic clk,
input logic reset,
input logic en,
input logic [WIDTH-1:0] d,
output logic [WIDTH-1:0] q
);
always_ff @(posedge clk or posedge reset)
if (reset) q <= {WIDTH{1'b0}};
else if (en) q <= d;
endmodule
